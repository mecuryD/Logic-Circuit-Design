module inv(input a,output z);

  assign z = ~a;
endmodule