module converter(rst,clk,data,ascii);

endmodule