module and1(a,b,z);
  input a;
  input b;
  output z;
  
  assign z = a&b;
endmodule